module
(

);






endmodule
